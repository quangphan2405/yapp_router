package yapp_pkg;

   import uvm_pkg::*;
`include "uvm_macros.svh"

`include "yapp_packet.sv"

endpackage : yapp_pkg
   
